`timescale 1ns / 1ps

module mux2 #(
    parameter WIDTH = 32
)(
    input [WIDTH-1:0] in0,  // Option 0
    input [WIDTH-1:0] in1,  // Option 1
    input sel, // Select line
    output [WIDTH-1:0]  out  // Output
);

assign out = (sel) ? in1 : in0;

endmodule
